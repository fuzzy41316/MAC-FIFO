module minilab1_2(
	//////////// CLOCK //////////
	input 		          		CLOCK2_50,
	input 		          		CLOCK3_50,
	input 		          		CLOCK4_50,
	input 		          		CLOCK_50,

	//////////// SEG7 //////////
	output	reg	     [6:0]		HEX0,
	output	reg	     [6:0]		HEX1,
	output	reg	     [6:0]		HEX2,
	output	reg	     [6:0]		HEX3,
	output	reg	     [6:0]		HEX4,
	output	reg	     [6:0]		HEX5,
	
	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// KEY //////////
	input 		     [3:0]		KEY,

	//////////// SW //////////
	input 		     [9:0]		SW
);
    

    // Internal wires
    /* SHARED */
    logic [7:0] datain;
    logic rst_n, Clr;

    /* MEMORY */
    reg [31:0] address;
    logic [63:0] readdata;
    logic readdatavalid, read;
    logic [7:0] readdata_byte [7:0];
    assign readdata_byte[0] = readdata[63:56];
    assign readdata_byte[1] = readdata[55:48];
    assign readdata_byte[2] = readdata[47:40];
    assign readdata_byte[3] = readdata[39:32];
    assign readdata_byte[4] = readdata[31:24];
    assign readdata_byte[5] = readdata[23:16];
    assign readdata_byte[6] = readdata[15:8];
    assign readdata_byte[7] = readdata[7:0];

    /* A ARRAY */
    logic [7:0] dataoutA [7:0];                 // Row of the 2D A array stored into the FIFO
    logic allFull;
    logic [7:0] rdenA, wrenA, emptyA, fullA;
    assign allFull = &fullA;

    /* B ARRAY */
    logic [7:0] dataoutB;                       // B array 
    logic rdenB, wrenB, emptyB, fullB;          // Control signals for the B FIFO

    /* MAC */
    logic [7:0] Ain;
    logic [7:0] Bin;
    logic [23:0] Cout [7:0];
    logic mac_count;    // TODO: increment the mac_count depending on the step you're on
                        // i.e., first Cout, then second Cout, then third Cout.
    
    // Instantiate the MAC module
    //TODO: tie inputs to mac directly to outputs from FIFO, control signals should come from SM
    mac mac(
        .clk(CLOCK_50),
        .rst_n(rst_n),
        .En(|rdenA & rdenB),    //TODO: Enable MAC if reading from B and any A?
        .Clr(Clr),
        .Ain(dataoutA[column]), //TODO:
        .Bin(dataoutB),         //TODO:
        .Cout(Cout[column]      //TODO: look here
        ));

    // Instantiate the memory module
    mem_wrapper memory(
        .clk(CLOCK_50),    
        .reset_n(rst_n),
        .address(address),              // 32-bit address for 8 rows
        .read(read),                    // Read request
        // Outputs
        .readdata(readdata),            // 64-bit read data (one row)
        .readdatavalid(readdatavalid),  // Data valid signal
        .waitrequest()                  // Busy signal to indicate logic is processing
    );


    // Generate FIFOs for the 8x8 A input
    genvar k;
    generate
    for (k = 0; k < 8; k++)  
    begin
        fifo A_fifo(
            .data(datain),
            .rdclk(CLOCK_50),
            .rdreq(rdenA[k]),
            .wrclk(CLOCK_50),
            .wrreq(wrenA[k]),
            // Outputs
            .q(dataoutA[k]),
            .rdempty(emptyA[k]),
            .wrfull(fullA[k])
        );
    end
    endgenerate

    generate
        begin
            fifo B_fifo(
                // Inputs
                .data(datain),
                .rdclk(CLOCK_50),
                .rdreq(rdenB),
                .wrclk(CLOCK_50),
                .wrreq(wrenB),
                // Outputs
                .q(dataoutB),
                .rdempty(emptyB),
                .wrfull(fullB)
            );
        end
    endgenerate

    // State and next state logic
    typedef enum reg [2:0] {READ, FILLA, FILLB, EXEC, DONE} state_t;
    state_t state, next_state;

    always_ff @(posedge CLOCK_50, negedge rst_n) 
    begin
        if (!rst_n)
            state <= READ;
        else 
            state <= next_state;
    end
    
    // Structural coding
    assign rst_n = KEY[0];
    logic reading;  // var to tell the column to start incrementing
    logic nextrow;  // For filling A

    // Counter for incrementing which byte-size column we're writing to the FIFO
    reg [2:0] column;
    always_ff@(posedge CLOCK_50, negedge rst_n) begin
        if (!rst_n) 
            column <= '0;
        else if (nextrow)
            column <= '0;
        else if (reading) 
            column <= column + 1;
        else if (fullB) 
            column <= '0;
    end

    // Counter for incrementing which byte-size column we're reading from the FIFO
    reg [2:0] row;
    always_ff@(posedge CLOCK_50, negedge rst_n) begin
        if (!rst_n) 
            row <= '0;
        else if (row_rst)
            row <= '0;
        else if (mac_exec) 
            row <= row + 1;
        else if (fullB) 
            row <= '0;
    end

    // ff to reset controlling signals on READ so we can reuse FILLB for mac
    //TODO: might have error with driving in two places in EXEC stage of SM
    reg mac_exec;
    always_ff@(posedge CLOCK_50, negedge rst_n) begin 
        if (!rst_n)
            mac_exec <= '0;
    end

    // Counter for address, to increment rows
    always_ff @(posedge CLOCK_50, negedge rst_n) begin
        if (!rst_n)
            address <= '0;
        else if (nextrow)
            address <= address + 1;
    end

    // State machine
    always_comb
    begin
        // Defaults
        read = '0;
        next_state = state;
        reading = 0;
        nextrow = 0;

        if (!rst_n)
        begin
            // Reset the FIFOs, start filling B first
            datain = '0;
            next_state = READ;
            wrenB = 0;
            rdenB = 0;
            wrenA = '0;
            rdenA = '0;
        end

        case(state)
            READ:
            begin
                read = 1'b1;
                // Need to check for data_valid signal from memory before filling the FIFO               
                else if (readdatavalid & !fullB)        // Fill B first
                    next_state = FILLB;
                else if (readdatavalid & !(allFull))    // Fill A second
                    next_state = FILLA;
                else if (fullB & allFull) begin         // Can start MAC
                    row_rst = '1;                       // assertion to reset the row counter after 
                    next_state = EXEC;
                end
            end

            FILLB:
            begin
                // As long as B FIFO is not full, keep filling
                if (!fullB) begin
                    reading = 1;
                    wrenB = 1'b1;
                    datain = readdata_byte[column];
                end
                else if (mac_exec) 
                    next_state = EXEC;   
                else begin
                    next_state = READ;
                    nextrow = 1;
                end
            end
            FILLA:
            begin
                if(!allFull)
                begin
                    reading = 1;
                    wrenA |= (1 << (address-1));
                    datain = readdata_byte[column];

                    // Read the next row
                    if (column == 7)
                    begin
                        nextrow = 1; 
                        wrenA |= (1 << (address-1));    
                        next_state = READ;
                    end
                end
            end
            
            EXEC:
            begin
                mac_exec = '1;
                // assert read signals;
                rdenA = '1;
                rdenB = '1;

                /*  NOTE: this is me exploiting the logic we already have here. will need other logic to support 
                    the interface between mac completing one entry in A (the 8 cycles it will take to read) and 
                    incrementing the counter to indicate which column we need to read from

                    by the time we get here, the logic for filling A is no longer needed. I want to reuse it to 
                    count where we are within each colcumn for reading. 
                */

                // logic to put the output of B FIFO into a 64 bit array so fill B can readd it to the FIFO
                readdata = readdata << 8;
                readdata |= dataoutB;
                if (&row) begin   //row == 7
                    
                    next_state = FILLB;
                end

            end
            
            DONE: 
            begin 
                // TODO: 
            end
            
            default:
            begin end 

        endcase
    end
endmodule