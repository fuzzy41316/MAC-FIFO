module testbench();




endmodule